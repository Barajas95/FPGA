LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SYNC IS
	PORT(	CLK: IN STD_LOGIC;
			HSYNC: OUT STD_LOGIC;
			VSYNC: OUT STD_LOGIC;
			R: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			G: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			B: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END SYNC;

ARCHITECTURE MAIN OF SYNC IS
	SIGNAL HPOS: INTEGER RANGE 0 TO 800:=0;
	SIGNAL VPOS: INTEGER RANGE 0 TO 525:=0;
BEGIN

PROCESS(CLK)
BEGIN
	IF(CLK'EVENT AND CLK='1') THEN
	
---------------------------------

		IF((VPOS>44 AND VPOS<141) OR (VPOS>237 AND VPOS<333) OR (VPOS>429 AND VPOS<525)) THEN
			R<="0000000000";		-- AZUL
			G<="0010101000";
			B<="1000111110";
		ELSE
			R<="1111111111";		-- BLANCO
			G<="1111111111";
			B<="1111111111";
		END IF;

		IF((HPOS-120)<VPOS AND VPOS<286) THEN
			R<="1100111110";		--ROJO
			G<="0001010000";
			B<="0010101100";
		END IF;
		
		IF(VPOS+HPOS<690 AND VPOS>285 AND HPOS<480) THEN
			R<="1100111110";		--ROJO
			G<="0001010000";
			B<="0010101100";
		END IF;
------		
		IF((VPOS=240 OR VPOS=239 OR VPOS=238) AND HPOS>251 AND HPOS<253) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=243 OR VPOS=242 OR VPOS=241) AND HPOS>250 AND HPOS<254) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=246 OR VPOS=245 OR VPOS=244) AND HPOS>249 AND HPOS<255) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=249 OR VPOS=248 OR VPOS=247) AND HPOS>248 AND HPOS<256) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=252 OR VPOS=251 OR VPOS=250) AND HPOS>247 AND HPOS<257) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=255 OR VPOS=254 OR VPOS=253) AND HPOS>246 AND HPOS<258) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=258 OR VPOS=257 OR VPOS=256) AND HPOS>245 AND HPOS<259) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=261 OR VPOS=260 OR VPOS=259) AND HPOS>244 AND HPOS<260) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=264 OR VPOS=263 OR VPOS=262) AND HPOS>243 AND HPOS<261) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=267 OR VPOS=266 OR VPOS=265) AND HPOS>242 AND HPOS<262) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=270 OR VPOS=269 OR VPOS=268) AND HPOS>241 AND HPOS<263) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
------
		IF(VPOS=271 AND HPOS>210 AND HPOS<294) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=272 AND HPOS>211 AND HPOS<293) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=273 AND HPOS>212 AND HPOS<292) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=274 AND HPOS>213 AND HPOS<291) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=275 AND HPOS>214 AND HPOS<290) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=276 AND HPOS>215 AND HPOS<289) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=277 AND HPOS>216 AND HPOS<288) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=278 AND HPOS>217 AND HPOS<287) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=279 AND HPOS>218 AND HPOS<286) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=280 AND HPOS>219 AND HPOS<285) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=281 AND HPOS>220 AND HPOS<284) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=282 AND HPOS>221 AND HPOS<283) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=283 AND HPOS>222 AND HPOS<282) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=284 AND HPOS>223 AND HPOS<281) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=285 AND HPOS>224 AND HPOS<280) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=286 AND HPOS>225 AND HPOS<279) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=287 AND HPOS>226 AND HPOS<278) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=288 AND HPOS>227 AND HPOS<277) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=289 AND HPOS>228 AND HPOS<276) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=290 AND HPOS>229 AND HPOS<275) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=291 AND HPOS>231 AND HPOS<274) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=292 AND HPOS>232 AND HPOS<273) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=293 AND HPOS>233 AND HPOS<272) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=294 AND HPOS>234 AND HPOS<271) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF(VPOS=295 AND HPOS>235 AND HPOS<270) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
------
		IF((VPOS=296 OR VPOS=297 OR VPOS=298) AND HPOS>234 AND HPOS<271) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=299 OR VPOS=300 OR VPOS=301) AND HPOS>233 AND HPOS<272) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=302 OR VPOS=303 OR VPOS=304) AND HPOS>232 AND HPOS<273) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=305 OR VPOS=306 OR VPOS=307) AND HPOS>231 AND HPOS<274) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=308 OR VPOS=309 OR VPOS=310) AND HPOS>230 AND HPOS<275) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
------
		IF((VPOS=311 OR VPOS=312 OR VPOS=313) AND ((HPOS>229 AND HPOS<251) OR (HPOS>252 AND HPOS<276))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=314 OR VPOS=315 OR VPOS=316) AND ((HPOS>228 AND HPOS<247) OR (HPOS>256 AND HPOS<277))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=317 OR VPOS=318 OR VPOS=319) AND ((HPOS>227 AND HPOS<243) OR (HPOS>260 AND HPOS<278))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=320 OR VPOS=321 OR VPOS=322) AND ((HPOS>226 AND HPOS<239) OR (HPOS>264 AND HPOS<279))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=323 OR VPOS=324 OR VPOS=325) AND ((HPOS>225 AND HPOS<235) OR (HPOS>268 AND HPOS<280))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=326 OR VPOS=327 OR VPOS=328) AND ((HPOS>224 AND HPOS<231) OR (HPOS>272 AND HPOS<281))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=329 OR VPOS=330 OR VPOS=331) AND ((HPOS>223 AND HPOS<227) OR (HPOS>276 AND HPOS<282))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=332 OR VPOS=333 OR VPOS=334) AND ((HPOS>222 AND HPOS<223) OR (HPOS>280 AND HPOS<283))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=335 OR VPOS=336 OR VPOS=337) AND ((HPOS>221 AND HPOS<219) OR (HPOS>284 AND HPOS<284))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		IF((VPOS=338 OR VPOS=339 OR VPOS=340) AND ((HPOS>220 AND HPOS<215) OR (HPOS>288 AND HPOS<285))) THEN
			R<="1111111111"; G<="1111111111"; B<="1111111111";
		END IF;
		
-------------------------------

		IF (HPOS<800) THEN
			HPOS<=HPOS+1;
		ELSE
			HPOS<=0;
			IF (VPOS<525) THEN
				VPOS<=VPOS+1;
			ELSE
				VPOS<=0;
			END IF;
		END IF;
	END IF;
	
---------------------------------

	IF(HPOS>16 AND HPOS<112) THEN
		HSYNC<='0';
	ELSE
		HSYNC<='1';
	END IF;
	
	IF(VPOS>10 AND VPOS<12) THEN
		VSYNC<='0';
	ELSE
		VSYNC<='1';
	END IF;
	
	IF((HPOS>0 AND HPOS<160) OR (VPOS>0 AND VPOS<45)) THEN		--PINTAR NEGRO EN LOS RANGOS FUERA DE LA PANTALLA
		R<="0000000000";
		G<="0000000000";
		B<="0000000000";
	END IF;
	
END PROCESS;

END MAIN;