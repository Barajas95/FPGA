LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FRECUENCIA4HZ IS
PORT(CLKIN: IN STD_LOGIC;
     CLKOUT: OUT STD_LOGIC);
END FRECUENCIA4HZ;

ARCHITECTURE RTL OF FRECUENCIA4HZ IS
	SIGNAL CICLOS: INTEGER RANGE 0 TO 6250000:=0;
BEGIN

PROCESS(CLKIN)
BEGIN
	IF(CLKIN'EVENT AND CLKIN = '1') THEN
		IF(CICLOS < 3125000) THEN
			CLKOUT <= '0';
			CICLOS<= CICLOS + 1;
		ELSE
			CLKOUT <= '1';
			CICLOS<= CICLOS + 1;
			IF(CICLOS=6250000)THEN
				CICLOS<=0;
			END IF;
		END IF;
	END IF;
END PROCESS;
END RTL;
