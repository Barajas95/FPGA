LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIVISOR_FRECUENCIA IS
PORT(CLKIN: IN STD_LOGIC;
     CLKOUT: OUT STD_LOGIC);
END DIVISOR_FRECUENCIA;

ARCHITECTURE RTL OF DIVISOR_FRECUENCIA IS
	SIGNAL CICLOS: INTEGER RANGE 0 TO 1:=0;
BEGIN

PROCESS(CLKIN)
BEGIN
	IF(CLKIN'EVENT AND CLKIN = '1') THEN
		IF(CICLOS = 0) THEN
			CLKOUT <= '0';
			CICLOS <= 1;
		ELSE
			CLKOUT <= '1';
			CICLOS<=0;
		END IF;
	END IF;
END PROCESS;
END RTL;
