LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY VGA IS
	PORT(	CLOCK_50: IN STD_LOGIC;
			VGA_HS: OUT STD_LOGIC;
			VGA_VS: OUT STD_LOGIC;
			VGA_R: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			VGA_G: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			VGA_B: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			BLANK: OUT STD_LOGIC;
			SINC: OUT STD_LOGIC;
			CLOCK_25: OUT STD_LOGIC);
END VGA;

ARCHITECTURE MAIN OF VGA IS
	
	SIGNAL VGACLK: STD_LOGIC;
	
	COMPONENT SYNC IS
		PORT(	CLK: IN STD_LOGIC;
				HSYNC: OUT STD_LOGIC;
				VSYNC: OUT STD_LOGIC;
				R: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
				G: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
				B: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
	END COMPONENT SYNC;
	
	COMPONENT DIVISOR_FRECUENCIA IS
		PORT(	CLKIN: IN STD_LOGIC;
				CLKOUT: OUT STD_LOGIC); 
	END COMPONENT DIVISOR_FRECUENCIA;
	
BEGIN
	C1: DIVISOR_FRECUENCIA PORT MAP(CLOCK_50,VGACLK);
	C2: SYNC PORT MAP(VGACLK,VGA_HS,VGA_VS,VGA_R,VGA_G,VGA_B);
	
	CLOCK_25<=VGACLK;
	BLANK<='1';
	SINC<='0';
	
END MAIN;