library verilog;
use verilog.vl_types.all;
entity Restador1_vlg_vec_tst is
end Restador1_vlg_vec_tst;
