LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY VGA IS
	PORT(	CLOCK_50: IN STD_LOGIC;
			PUSH_YELLOW: IN STD_LOGIC;
			PUSH_BLUE: IN STD_LOGIC;
			PUSH_RED: IN STD_LOGIC;
			PUSH_GREEN: IN STD_LOGIC;
			SWITCH_PRENDIDOAPAGADO: IN STD_LOGIC;
			SWITCH_NIVEL1: IN STD_LOGIC;
			SWITCH_NIVEL2: IN STD_LOGIC;
			SWITCH_NIVEL3: IN STD_LOGIC;
			VGA_HS: OUT STD_LOGIC;
			VGA_VS: OUT STD_LOGIC;
			VGA_R: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			VGA_G: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			VGA_B: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			BLANK: OUT STD_LOGIC;
			SINC: OUT STD_LOGIC;
			CLOCK_25: OUT STD_LOGIC);
END VGA;

ARCHITECTURE MAIN OF VGA IS
	
	SIGNAL VGACLK25: STD_LOGIC;
	SIGNAL VGACLK2HZ: STD_LOGIC;
	SIGNAL VGACLK4HZ: STD_LOGIC;
	SIGNAL VGACLK8HZ: STD_LOGIC;
	SIGNAL VELOCIDAD: STD_LOGIC;
	SIGNAL VGAPOSICIONH: INTEGER RANGE 0 TO 800:=0;
	SIGNAL VGAPOSICIONV: INTEGER RANGE 0 TO 525:=0;
	
	COMPONENT SYNC IS
		PORT(	CLK: IN STD_LOGIC;
				HSYNC: OUT STD_LOGIC;
				VSYNC: OUT STD_LOGIC;
				VALORH: OUT INTEGER RANGE 0 TO 800;
				VALORV: OUT INTEGER RANGE 0 TO 525);
	END COMPONENT SYNC;
	
	COMPONENT DIVISOR_FRECUENCIA IS
		PORT(	CLKIN: IN STD_LOGIC;
				CLKOUT: OUT STD_LOGIC); 
	END COMPONENT DIVISOR_FRECUENCIA;
	
	COMPONENT FRECUENCIA2HZ IS
		PORT(	CLKIN: IN STD_LOGIC;
				CLKOUT: OUT STD_LOGIC); 
	END COMPONENT FRECUENCIA2HZ;
	
	COMPONENT FRECUENCIA4HZ IS
		PORT(	CLKIN: IN STD_LOGIC;
				CLKOUT: OUT STD_LOGIC); 
	END COMPONENT FRECUENCIA4HZ;

	COMPONENT FRECUENCIA8HZ IS
		PORT(	CLKIN: IN STD_LOGIC;
				CLKOUT: OUT STD_LOGIC); 
	END COMPONENT FRECUENCIA8HZ;
	
	COMPONENT MULTIPLEXORSIMON IS
		PORT(	CLK1: IN STD_LOGIC;
				CLK2: IN STD_LOGIC;
				CLK3: IN STD_LOGIC;
				PUSH1: IN STD_LOGIC;
				PUSH2: IN STD_LOGIC;
				PUSH3: IN STD_LOGIC;
				PUSH_ONOFF: IN STD_LOGIC;
				SALIDA: OUT STD_LOGIC);
	END COMPONENT MULTIPLEXORSIMON;
	
	COMPONENT PANTALLA IS
		PORT(	VALORH: IN INTEGER RANGE 0 TO 800;
				VALORV: IN INTEGER RANGE 0 TO 525;
				PUSH_AMARILLO: IN STD_LOGIC;
				PUSH_AZUL: IN STD_LOGIC;
				PUSH_ROJO: IN STD_LOGIC;
				PUSH_VERDE: IN STD_LOGIC;
				SWITCH_ONOFF: IN STD_LOGIC;
				SWITCH_LEVEL1: IN STD_LOGIC;
				SWITCH_LEVEL2: IN STD_LOGIC;
				SWITCH_LEVEL3: IN STD_LOGIC;
				CLOCK25MHZ: IN STD_LOGIC;
				VELOCIDAD: IN STD_LOGIC;
				R: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
				G: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
				B: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
	END COMPONENT PANTALLA;
BEGIN
	D1: DIVISOR_FRECUENCIA PORT MAP(CLOCK_50,VGACLK25);
	D2: FRECUENCIA2HZ PORT MAP(VGACLK25,VGACLK2HZ);
	D3: FRECUENCIA4HZ PORT MAP (VGACLK25,VGACLK4HZ);
	D4: FRECUENCIA8HZ PORT MAP (VGACLK25,VGACLK8HZ);
	D5: MULTIPLEXORSIMON PORT MAP(VGACLK2HZ,VGACLK4HZ,VGACLK8HZ,SWITCH_NIVEL1,SWITCH_NIVEL2,SWITCH_NIVEL3,SWITCH_PRENDIDOAPAGADO,VELOCIDAD);
	
	C1: SYNC PORT MAP(VGACLK25,VGA_HS,VGA_VS,VGAPOSICIONH,VGAPOSICIONV);
	C2: PANTALLA PORT MAP(VGAPOSICIONH,VGAPOSICIONV,PUSH_YELLOW,PUSH_BLUE,PUSH_RED,PUSH_GREEN,SWITCH_PRENDIDOAPAGADO,SWITCH_NIVEL1,SWITCH_NIVEL2,SWITCH_NIVEL3,VGACLK25,VELOCIDAD,VGA_R,VGA_G,VGA_B);
	
	CLOCK_25<=VGACLK25;
	BLANK<='1';
	SINC<='0';
	
END MAIN;