library verilog;
use verilog.vl_types.all;
entity VGA_vlg_vec_tst is
end VGA_vlg_vec_tst;
