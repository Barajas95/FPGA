LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SYNC IS
	PORT(	CLK: IN STD_LOGIC;
			HSYNC: OUT STD_LOGIC;
			VSYNC: OUT STD_LOGIC;
			VALORH: OUT INTEGER RANGE 0 TO 800;
			VALORV: OUT INTEGER RANGE 0 TO 525);
END SYNC;

ARCHITECTURE MAIN OF SYNC IS
	SIGNAL HPOS: INTEGER RANGE 0 TO 800:=0;
	SIGNAL VPOS: INTEGER RANGE 0 TO 525:=0;
BEGIN

PROCESS(CLK)
BEGIN
	IF(CLK'EVENT AND CLK='1') THEN
		IF (HPOS<800) THEN
			HPOS<=HPOS+1;
		ELSE
			HPOS<=0;
			IF (VPOS<525) THEN
				VPOS<=VPOS+1;
			ELSE
				VPOS<=0;
			END IF;
		END IF;		
	END IF;

	IF(HPOS>16 AND HPOS<112) THEN
		HSYNC<='0';
	ELSE
		HSYNC<='1';
	END IF;
	
	IF(VPOS>10 AND VPOS<12) THEN
		VSYNC<='0';
	ELSE
		VSYNC<='1';
	END IF;
	
	VALORH<=HPOS;
	VALORV<=VPOS;
	
END PROCESS;

END MAIN;